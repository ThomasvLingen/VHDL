----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:52:21 03/11/2015 
-- Design Name: 
-- Module Name:    soundByteSelector - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity soundByteSelector is
    Port ( sampleCounter : in  STD_LOGIC_VECTOR(11 downto 0);
			  clk25 : in STD_LOGIC;
           soundByte : out  STD_LOGIC_VECTOR(7 downto 0));
end soundByteSelector;

architecture Behavioral of soundByteSelector is

begin

	process(clk25, sampleCounter)
		variable currentByte : integer := 0;
		type RomType is array (natural range <>) of std_logic_vector(7 downto 0);
		
		constant soundLength: integer := 6667;
		
		constant Sound: RomType(0 to 6667) := (
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"81", X"81", X"80", X"80", X"80", X"80", X"80", X"81", X"81", X"80", X"80", X"80", X"80", 
		X"80", X"81", X"80", X"81", X"80", X"80", X"81", X"80", X"80", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"81", X"81", X"81", X"81", X"81", X"80", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"81", X"81", X"80", 
		X"80", X"80", X"80", X"80", X"81", X"81", X"80", X"81", X"80", X"80", X"80", X"80", X"81", X"80", X"81", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"81", X"80", X"81", X"80", X"7f", X"7f", X"7f", X"80", X"80", X"80", 
		X"80", X"7f", X"7f", X"7f", X"7f", X"80", X"80", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7e", X"7f", 
		X"7f", X"7f", X"80", X"7f", X"7e", X"7d", X"7d", X"7d", X"7e", X"7f", X"7f", X"80", X"80", X"7f", X"7e", X"7d", 
		X"7c", X"7c", X"7f", X"81", X"83", X"83", X"81", X"7f", X"7e", X"7f", X"7f", X"80", X"81", X"82", X"83", X"83", 
		X"83", X"83", X"82", X"81", X"81", X"82", X"82", X"83", X"83", X"83", X"83", X"83", X"82", X"81", X"81", X"81", 
		X"82", X"82", X"83", X"82", X"82", X"82", X"81", X"81", X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"80", 
		X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7e", X"7e", X"7d", X"7c", X"7c", X"7c", X"7b", X"7b", X"7b", X"7b", 
		X"7c", X"7d", X"7e", X"7e", X"7d", X"7d", X"7d", X"7f", X"81", X"81", X"80", X"7e", X"7f", X"81", X"84", X"85", 
		X"84", X"84", X"82", X"82", X"84", X"84", X"85", X"84", X"85", X"86", X"86", X"86", X"86", X"85", X"85", X"84", 
		X"85", X"85", X"84", X"84", X"84", X"83", X"83", X"83", X"83", X"83", X"82", X"81", X"80", X"7f", X"80", X"7f", 
		X"7e", X"7f", X"7e", X"7e", X"7d", X"7d", X"7d", X"7c", X"7b", X"79", X"77", X"78", X"76", X"77", X"79", X"7a", 
		X"7d", X"7e", X"7e", X"7d", X"7b", X"79", X"79", X"7a", X"7b", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"80", X"80", X"81", X"83", X"83", X"84", X"85", X"85", X"85", X"85", X"85", X"84", X"85", X"86", X"86", X"87", 
		X"86", X"86", X"85", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"83", X"82", X"81", X"81", X"7f", X"7e", 
		X"7e", X"7d", X"7d", X"7d", X"7c", X"7c", X"79", X"79", X"77", X"75", X"78", X"78", X"7e", X"7f", X"80", X"7f", 
		X"7b", X"7b", X"78", X"78", X"79", X"7b", X"7e", X"7f", X"81", X"81", X"81", X"7f", X"7e", X"7d", X"7d", X"7f", 
		X"82", X"84", X"87", X"88", X"87", X"87", X"86", X"85", X"84", X"85", X"86", X"87", X"89", X"89", X"89", X"88", 
		X"86", X"84", X"84", X"84", X"85", X"86", X"86", X"85", X"83", X"81", X"80", X"7e", X"7d", X"7c", X"7c", X"7c", 
		X"7d", X"7c", X"78", X"75", X"71", X"78", X"7f", X"85", X"8a", X"84", X"7e", X"77", X"75", X"75", X"78", X"7b", 
		X"7b", X"7d", X"7f", X"80", X"83", X"83", X"82", X"7d", X"7c", X"7a", X"7b", X"80", X"83", X"87", X"87", X"87", 
		X"86", X"85", X"85", X"85", X"85", X"85", X"85", X"85", X"86", X"86", X"86", X"84", X"82", X"81", X"81", X"82", 
		X"82", X"81", X"7f", X"7c", X"7c", X"7b", X"7a", X"79", X"77", X"73", X"71", X"75", X"7b", X"88", X"8b", X"8a", 
		X"84", X"78", X"74", X"71", X"75", X"79", X"7c", X"80", X"81", X"84", X"86", X"85", X"83", X"7d", X"79", X"77", 
		X"77", X"7a", X"81", X"87", X"8a", X"8d", X"8a", X"88", X"85", X"82", X"81", X"81", X"82", X"84", X"88", X"8a", 
		X"89", X"87", X"82", X"7e", X"7c", X"7d", X"7f", X"80", X"81", X"7e", X"7c", X"78", X"75", X"74", X"6e", X"6c", 
		X"73", X"82", X"8d", X"94", X"90", X"82", X"76", X"70", X"6e", X"73", X"79", X"7d", X"81", X"86", X"8a", X"8c", 
		X"8d", X"87", X"7e", X"76", X"73", X"74", X"78", X"81", X"8a", X"91", X"96", X"93", X"8e", X"86", X"80", X"7d", 
		X"7e", X"83", X"87", X"8d", X"8f", X"8d", X"89", X"83", X"7e", X"7d", X"7e", X"7f", X"7f", X"7c", X"78", X"73", 
		X"71", X"71", X"70", X"76", X"88", X"8d", X"90", X"8f", X"7f", X"77", X"6f", X"6e", X"6e", X"73", X"79", X"7c", 
		X"87", X"8f", X"91", X"8f", X"84", X"76", X"6d", X"6b", X"6f", X"79", X"86", X"8f", X"97", X"97", X"91", X"89", 
		X"7f", X"7a", X"79", X"7d", X"84", X"8b", X"8f", X"90", X"8c", X"85", X"7f", X"7b", X"79", X"7b", X"7d", X"7b", 
		X"76", X"71", X"6d", X"69", X"7b", X"95", X"92", X"9a", X"89", X"74", X"70", X"6e", X"75", X"74", X"7b", X"78", 
		X"78", X"85", X"88", X"8d", X"8f", X"82", X"75", X"6e", X"6b", X"70", X"7d", X"8a", X"8f", X"93", X"8e", X"87", 
		X"83", X"7f", X"7d", X"7d", X"7e", X"81", X"86", X"8a", X"88", X"83", X"7c", X"77", X"77", X"7b", X"7a", X"78", 
		X"74", X"6a", X"66", X"80", X"96", X"94", X"a3", X"85", X"73", X"6f", X"6c", X"7a", X"7c", X"87", X"7c", X"7c", 
		X"86", X"84", X"92", X"90", X"83", X"79", X"71", X"6f", X"77", X"89", X"90", X"95", X"93", X"87", X"82", X"80", 
		X"80", X"81", X"84", X"83", X"83", X"87", X"84", X"80", X"79", X"72", X"6d", X"6f", X"76", X"79", X"77", X"75", 
		X"7f", X"8b", X"8c", X"93", X"7e", X"72", X"6a", X"69", X"78", X"80", X"8c", X"88", X"86", X"84", X"7f", X"85", 
		X"82", X"7e", X"7a", X"77", X"7b", X"86", X"91", X"97", X"96", X"8d", X"83", X"7d", X"7e", X"83", X"88", X"8c", 
		X"8c", X"8a", X"87", X"80", X"7a", X"74", X"70", X"70", X"6f", X"6d", X"6c", X"77", X"98", X"98", X"9f", X"95", 
		X"6a", X"6a", X"59", X"69", X"74", X"7f", X"87", X"7c", X"8c", X"84", X"8b", X"8d", X"7b", X"71", X"67", X"6a", 
		X"75", X"8c", X"96", X"98", X"94", X"84", X"7e", X"7b", X"7d", X"7f", X"84", X"84", X"85", X"88", X"82", X"7c", 
		X"72", X"6c", X"68", X"68", X"6a", X"78", X"9b", X"9d", X"a4", X"9a", X"71", X"6c", X"57", X"65", X"6d", X"7d", 
		X"89", X"85", X"96", X"90", X"94", X"8f", X"7b", X"6e", X"64", X"67", X"73", X"8a", X"97", X"9d", X"9a", X"8a", 
		X"80", X"77", X"76", X"77", X"7d", X"82", X"86", X"87", X"80", X"76", X"6c", X"67", X"65", X"65", X"6e", X"89", 
		X"9b", X"9d", X"a1", X"81", X"70", X"63", X"5f", X"6b", X"72", X"83", X"82", X"8f", X"93", X"92", X"95", X"85", 
		X"76", X"69", X"69", X"72", X"86", X"96", X"9d", X"9e", X"91", X"86", X"7e", X"7a", X"7a", X"7f", X"84", X"86", 
		X"88", X"80", X"77", X"6f", X"6a", X"65", X"69", X"7a", X"91", X"99", X"a0", X"91", X"77", X"6e", X"5f", X"65", 
		X"6c", X"76", X"7f", X"86", X"91", X"91", X"95", X"8d", X"7c", X"70", X"66", X"6b", X"77", X"89", X"95", X"9b", 
		X"98", X"8d", X"83", X"7a", X"76", X"77", X"7c", X"80", X"85", X"82", X"7a", X"71", X"6c", X"67", X"6a", X"7b", 
		X"92", X"98", X"9c", X"91", X"76", X"6e", X"63", X"67", X"6d", X"75", X"7d", X"82", X"90", X"91", X"96", X"8f", 
		X"7e", X"6f", X"66", X"69", X"76", X"8a", X"93", X"9a", X"96", X"8d", X"84", X"7d", X"78", X"77", X"7a", X"7c", 
		X"7f", X"7d", X"74", X"6d", X"69", X"65", X"70", X"86", X"94", X"99", X"96", X"81", X"6f", X"67", X"62", X"68", 
		X"6f", X"76", X"7d", X"88", X"91", X"95", X"94", X"88", X"77", X"6a", X"66", X"6d", X"7d", X"8c", X"95", X"99", 
		X"94", X"8b", X"84", X"7d", X"79", X"79", X"7b", X"7e", X"7e", X"79", X"70", X"6c", X"6a", X"6c", X"82", X"95", 
		X"9a", X"9c", X"8a", X"72", X"69", X"61", X"67", X"6e", X"75", X"7b", X"83", X"8f", X"94", X"98", X"8f", X"7e", 
		X"6e", X"65", X"69", X"78", X"8a", X"93", X"98", X"94", X"8c", X"86", X"80", X"7c", X"7b", X"7c", X"7d", X"7d", 
		X"79", X"71", X"6d", X"6b", X"6d", X"80", X"98", X"9c", X"9f", X"90", X"74", X"6c", X"61", X"65", X"6b", X"74", 
		X"7b", X"82", X"90", X"93", X"96", X"8f", X"7d", X"6e", X"66", X"68", X"75", X"87", X"90", X"96", X"92", X"8c", 
		X"86", X"80", X"7b", X"78", X"79", X"79", X"7c", X"78", X"71", X"6c", X"69", X"6b", X"7f", X"98", X"9d", X"a1", 
		X"8f", X"74", X"6b", X"62", X"67", X"6e", X"76", X"7b", X"83", X"90", X"94", X"98", X"90", X"7d", X"6e", X"66", 
		X"69", X"77", X"88", X"90", X"94", X"8f", X"87", X"82", X"7c", X"78", X"76", X"77", X"78", X"78", X"73", X"69", 
		X"65", X"61", X"66", X"84", X"99", X"9e", X"a2", X"87", X"6f", X"65", X"5d", X"65", X"6c", X"77", X"7a", X"87", 
		X"94", X"98", X"9c", X"8e", X"79", X"69", X"62", X"68", X"7c", X"8d", X"96", X"9a", X"92", X"89", X"82", X"7d", 
		X"78", X"78", X"77", X"78", X"78", X"73", X"6b", X"66", X"62", X"6a", X"8a", X"98", X"9e", X"9d", X"7d", X"70", 
		X"63", X"61", X"67", X"6b", X"74", X"76", X"88", X"93", X"9b", X"9d", X"8b", X"77", X"67", X"63", X"6c", X"80", 
		X"8e", X"97", X"97", X"8f", X"89", X"83", X"7d", X"79", X"78", X"77", X"78", X"76", X"6f", X"69", X"66", X"65", 
		X"7c", X"97", X"99", X"a1", X"8d", X"72", X"6b", X"60", X"67", X"6a", X"72", X"75", X"7e", X"8f", X"95", X"9d", 
		X"95", X"82", X"6f", X"65", X"67", X"76", X"88", X"91", X"97", X"91", X"8a", X"85", X"80", X"7c", X"79", X"77", 
		X"76", X"77", X"72", X"6c", X"68", X"64", X"6b", X"8d", X"97", X"9f", X"9e", X"7c", X"6f", X"60", X"5f", X"66", 
		X"6d", X"74", X"76", X"86", X"8e", X"97", X"9a", X"8b", X"79", X"6a", X"64", X"6b", X"7e", X"8b", X"95", X"95", 
		X"8e", X"88", X"83", X"7d", X"79", X"78", X"76", X"76", X"74", X"6d", X"68", X"65", X"63", X"79", X"94", X"97", 
		X"a3", X"8d", X"74", X"6b", X"5e", X"64", X"66", X"70", X"72", X"7c", X"8a", X"91", X"9b", X"93", X"82", X"70", 
		X"66", X"66", X"74", X"86", X"91", X"98", X"92", X"8a", X"83", X"7f", X"7b", X"7a", X"79", X"77", X"77", X"73", 
		X"6d", X"67", X"63", X"6c", X"8b", X"94", X"9c", X"99", X"7c", X"73", X"67", X"67", X"69", X"6c", X"70", X"72", 
		X"82", X"8c", X"98", X"9a", X"8b", X"7a", X"6b", X"66", X"6d", X"7f", X"8b", X"95", X"95", X"8f", X"8a", X"85", 
		X"80", X"7c", X"7a", X"78", X"7a", X"79", X"73", X"6d", X"68", X"64", X"73", X"90", X"97", X"a2", X"96", X"7a", 
		X"70", X"63", X"66", X"69", X"70", X"72", X"77", X"87", X"8f", X"9b", X"9a", X"8a", X"78", X"68", X"63", X"6e", 
		X"81", X"8e", X"99", X"97", X"90", X"89", X"83", X"7d", X"79", X"77", X"75", X"77", X"74", X"6f", X"6b", X"68", 
		X"72", X"90", X"97", X"9c", X"97", X"79", X"72", X"69", X"6b", X"6e", X"70", X"72", X"71", X"81", X"8a", X"97", 
		X"9b", X"8d", X"7c", X"6e", X"68", X"6d", X"7e", X"88", X"91", X"92", X"8d", X"8b", X"87", X"82", X"7c", X"79", 
		X"75", X"75", X"73", X"6d", X"68", X"65", X"6c", X"89", X"98", X"9e", X"9e", X"82", X"74", X"68", X"66", X"69", 
		X"6c", X"71", X"70", X"7f", X"8a", X"96", X"9e", X"94", X"81", X"70", X"65", X"67", X"77", X"84", X"90", X"94", 
		X"90", X"8d", X"88", X"83", X"7c", X"78", X"73", X"73", X"72", X"6e", X"69", X"67", X"70", X"8c", X"99", X"9f", 
		X"9a", X"7f", X"73", X"6a", X"6b", X"6e", X"6f", X"70", X"6d", X"7b", X"87", X"96", X"9e", X"96", X"85", X"74", 
		X"6a", X"6b", X"79", X"83", X"8c", X"8f", X"8d", X"8d", X"8b", X"87", X"7f", X"79", X"74", X"71", X"6f", X"69", 
		X"65", X"66", X"77", X"93", X"9e", X"a5", X"98", X"7e", X"72", X"68", X"6d", X"6e", X"72", X"71", X"72", X"80", 
		X"8b", X"9a", X"9e", X"93", X"82", X"73", X"6b", X"70", X"7d", X"86", X"8e", X"8f", X"8e", X"8d", X"8c", X"86", 
		X"7e", X"77", X"71", X"6f", X"6c", X"66", X"63", X"6a", X"85", X"98", X"a1", X"a2", X"89", X"78", X"6c", X"68", 
		X"6d", X"6f", X"72", X"6e", X"78", X"84", X"91", X"9d", X"99", X"8c", X"7c", X"70", X"6d", X"76", X"80", X"87", 
		X"8d", X"8c", X"8d", X"8e", X"8c", X"85", X"7d", X"74", X"6e", X"6b", X"66", X"61", X"65", X"7b", X"93", X"9e", 
		X"a5", X"94", X"7e", X"71", X"68", X"68", X"69", X"6d", X"6c", X"73", X"82", X"8e", X"9a", X"9c", X"8f", X"80", 
		X"73", X"6b", X"71", X"7b", X"82", X"89", X"8c", X"8c", X"8e", X"8d", X"87", X"7e", X"76", X"6f", X"6a", X"67", 
		X"61", X"63", X"76", X"8f", X"9b", X"a5", X"99", X"83", X"77", X"6b", X"69", X"68", X"69", X"68", X"6d", X"7d", 
		X"8b", X"9a", X"a0", X"96", X"87", X"79", X"6f", X"70", X"79", X"7f", X"85", X"89", X"8b", X"8f", X"91", X"8c", 
		X"83", X"78", X"6f", X"68", X"64", X"60", X"62", X"78", X"8f", X"9a", X"a5", X"9a", X"88", X"7d", X"72", X"6c", 
		X"68", X"67", X"63", X"6a", X"79", X"89", X"99", X"a1", X"99", X"8b", X"7f", X"73", X"71", X"77", X"7b", X"81", 
		X"86", X"8a", X"8e", X"93", X"8f", X"86", X"7d", X"71", X"68", X"62", X"5e", X"63", X"7b", X"8e", X"99", X"a3", 
		X"98", X"8b", X"82", X"78", X"6f", X"69", X"65", X"5f", X"67", X"76", X"85", X"96", X"9e", X"9a", X"91", X"86", 
		X"79", X"74", X"75", X"76", X"7b", X"82", X"88", X"8e", X"93", X"8f", X"88", X"7e", X"73", X"68", X"61", X"5e", 
		X"65", X"7b", X"8a", X"95", X"9c", X"94", X"8c", X"85", X"7d", X"74", X"6c", X"66", X"60", X"65", X"71", X"7d", 
		X"8c", X"95", X"95", X"92", X"8d", X"84", X"7d", X"79", X"74", X"75", X"7a", X"80", X"87", X"8d", X"8e", X"89", 
		X"82", X"79", X"6e", X"66", X"62", X"65", X"75", X"83", X"8c", X"95", X"91", X"8d", X"8a", X"84", X"7c", X"74", 
		X"6e", X"66", X"67", X"6e", X"75", X"80", X"89", X"8c", X"8e", X"8e", X"8b", X"86", X"83", X"7e", X"7b", X"7b", 
		X"7d", X"81", X"85", X"88", X"87", X"85", X"7f", X"76", X"6e", X"68", X"67", X"6e", X"7b", X"83", X"8a", X"8c", 
		X"8a", X"88", X"89", X"86", X"83", X"7e", X"76", X"6f", X"6f", X"71", X"75", X"7d", X"81", X"83", X"85", X"87", 
		X"88", X"8b", X"8d", X"8a", X"87", X"84", X"81", X"83", X"85", X"87", X"86", X"84", X"7e", X"77", X"71", X"6a", 
		X"68", X"6c", X"77", X"80", X"87", X"8c", X"8b", X"8a", X"8b", X"89", X"86", X"83", X"7c", X"76", X"72", X"72", 
		X"74", X"78", X"7d", X"7f", X"80", X"82", X"84", X"89", X"8e", X"8f", X"8e", X"8b", X"87", X"86", X"86", X"85", 
		X"84", X"81", X"7e", X"79", X"74", X"6d", X"6a", X"6b", X"72", X"7d", X"83", X"88", X"8a", X"89", X"89", X"8a", 
		X"89", X"86", X"82", X"7b", X"76", X"73", X"73", X"74", X"78", X"7b", X"7b", X"7e", X"80", X"84", X"8a", X"8e", 
		X"8f", X"8e", X"8c", X"88", X"86", X"85", X"83", X"81", X"7f", X"7c", X"77", X"71", X"6b", X"69", X"6c", X"75", 
		X"7d", X"82", X"86", X"87", X"86", X"88", X"89", X"88", X"87", X"82", X"7d", X"79", X"76", X"76", X"77", X"7a", 
		X"7a", X"7a", X"7b", X"7d", X"81", X"88", X"8d", X"90", X"90", X"8e", X"89", X"88", X"86", X"84", X"82", X"7f", 
		X"7a", X"76", X"72", X"6d", X"6b", X"6d", X"74", X"7b", X"7f", X"84", X"85", X"86", X"87", X"88", X"89", X"87", 
		X"85", X"81", X"7d", X"7b", X"7a", X"79", X"7a", X"7b", X"7a", X"7b", X"7e", X"82", X"88", X"8d", X"91", X"91", 
		X"90", X"8c", X"8a", X"89", X"87", X"84", X"81", X"7e", X"7a", X"77", X"72", X"6f", X"6e", X"71", X"78", X"7b", 
		X"81", X"84", X"85", X"87", X"87", X"89", X"88", X"88", X"86", X"82", X"7f", X"7b", X"7a", X"79", X"7a", X"7b", 
		X"7b", X"7d", X"7f", X"83", X"87", X"8c", X"8f", X"8f", X"8e", X"8b", X"89", X"88", X"86", X"85", X"83", X"80", 
		X"7c", X"77", X"72", X"6e", X"6e", X"73", X"78", X"7c", X"82", X"83", X"84", X"85", X"86", X"89", X"89", X"89", 
		X"87", X"83", X"80", X"7d", X"7c", X"7c", X"7c", X"7c", X"7c", X"7d", X"7e", X"81", X"85", X"88", X"8b", X"8c", 
		X"8b", X"89", X"89", X"89", X"87", X"86", X"83", X"7f", X"7c", X"77", X"72", X"6e", X"6c", X"6f", X"74", X"79", 
		X"7e", X"81", X"82", X"83", X"84", X"88", X"88", X"8a", X"89", X"85", X"82", X"7f", X"7d", X"7d", X"7d", X"7d", 
		X"7d", X"7d", X"7c", X"7e", X"80", X"84", X"88", X"8b", X"8d", X"8c", X"8b", X"8b", X"8a", X"89", X"88", X"84", 
		X"81", X"7b", X"76", X"70", X"6d", X"6e", X"72", X"77", X"7c", X"7f", X"80", X"82", X"83", X"86", X"89", X"89", 
		X"8a", X"87", X"85", X"82", X"80", X"81", X"80", X"80", X"7e", X"7b", X"7a", X"79", X"7b", X"80", X"85", X"8a", 
		X"8d", X"8e", X"8d", X"8c", X"8d", X"8c", X"8a", X"88", X"83", X"80", X"7d", X"79", X"76", X"72", X"70", X"73", 
		X"7a", X"7b", X"7f", X"83", X"83", X"86", X"88", X"8a", X"89", X"89", X"89", X"87", X"85", X"83", X"80", X"7e", 
		X"7d", X"7b", X"7c", X"7c", X"7c", X"7f", X"83", X"88", X"8d", X"90", X"90", X"8d", X"8b", X"89", X"87", X"88", 
		X"84", X"82", X"80", X"7c", X"77", X"71", X"6e", X"6c", X"73", X"81", X"86", X"8a", X"8d", X"88", X"8b", X"8b", 
		X"8a", X"88", X"83", X"7e", X"76", X"74", X"74", X"75", X"7a", X"7e", X"7e", X"82", X"85", X"8a", X"8e", X"92", 
		X"92", X"8d", X"8a", X"84", X"81", X"82", X"81", X"82", X"84", X"85", X"84", X"82", X"7f", X"78", X"72", X"6d", 
		X"6c", X"72", X"82", X"89", X"8d", X"92", X"89", X"8a", X"8a", X"88", X"85", X"7c", X"76", X"6b", X"6c", X"72", 
		X"77", X"82", X"87", X"87", X"89", X"8a", X"8d", X"8e", X"90", X"8a", X"81", X"7d", X"7a", X"7d", X"82", X"88", 
		X"8a", X"8c", X"8d", X"8c", X"8b", X"86", X"7f", X"77", X"71", X"6a", X"67", X"6a", X"75", X"84", X"8b", X"93", 
		X"92", X"8d", X"8e", X"8a", X"86", X"7e", X"76", X"6e", X"6b", X"71", X"77", X"7f", X"86", X"87", X"89", X"8b", 
		X"8e", X"90", X"90", X"8b", X"83", X"7e", X"7d", X"80", X"86", X"8b", X"8d", X"8c", X"8e", X"8d", X"8c", X"87", 
		X"7f", X"77", X"71", X"6c", X"68", X"69", X"73", X"83", X"8c", X"94", X"96", X"8e", X"8d", X"89", X"86", X"80", 
		X"78", X"71", X"6a", X"6e", X"75", X"7d", X"87", X"8a", X"8c", X"8d", X"8f", X"90", X"8f", X"8a", X"81", X"7a", 
		X"78", X"7b", X"83", X"8a", X"8e", X"8f", X"90", X"91", X"8e", X"8a", X"82", X"79", X"73", X"70", X"6c", X"68", 
		X"67", X"6e", X"7f", X"8d", X"97", X"9a", X"92", X"8d", X"87", X"84", X"7f", X"76", X"6f", X"66", X"68", X"72", 
		X"7d", X"8a", X"91", X"92", X"91", X"8f", X"8d", X"89", X"85", X"7c", X"74", X"73", X"78", X"81", X"8b", X"92", 
		X"93", X"93", X"92", X"8e", X"88", X"81", X"7a", X"74", X"73", X"70", X"6b", X"66", X"64", X"6b", X"7e", X"92", 
		X"99", X"9d", X"94", X"8a", X"85", X"82", X"7e", X"73", X"6b", X"63", X"63", X"72", X"81", X"8f", X"96", X"95", 
		X"8f", X"8a", X"89", X"86", X"81", X"7a", X"71", X"6e", X"75", X"81", X"8e", X"97", X"9a", X"96", X"91", X"8c", 
		X"87", X"81", X"7c", X"78", X"76", X"76", X"74", X"71", X"6d", X"6c", X"70", X"7f", X"92", X"98", X"99", X"94", 
		X"88", X"83", X"7f", X"7c", X"74", X"6c", X"68", X"68", X"75", X"85", X"91", X"97", X"95", X"8e", X"87", X"85", 
		X"83", X"7e", X"79", X"73", X"6e", X"74", X"82", X"8f", X"99", X"9d", X"99", X"92", X"8d", X"88", X"82", X"7e", 
		X"7b", X"79", X"7b", X"7c", X"77", X"73", X"6f", X"6d", X"72", X"7f", X"8f", X"94", X"94", X"92", X"86", X"82", 
		X"80", X"7c", X"75", X"6e", X"6d", X"6e", X"79", X"87", X"8e", X"92", X"90", X"88", X"83", X"81", X"80", X"7c", 
		X"7a", X"77", X"74", X"79", X"85", X"90", X"98", X"9c", X"98", X"8f", X"8a", X"84", X"7e", X"7b", X"7b", X"7a", 
		X"7c", X"7e", X"7a", X"75", X"71", X"6e", X"6d", X"73", X"80", X"8b", X"8e", X"91", X"8b", X"83", X"81", X"7d", 
		X"79", X"73", X"70", X"6e", X"70", X"7c", X"85", X"8c", X"8f", X"8c", X"86", X"83", X"81", X"7f", X"7c", X"7b", 
		X"78", X"77", X"7d", X"88", X"91", X"97", X"99", X"93", X"8b", X"86", X"80", X"7c", X"7b", X"7b", X"7b", X"7d", 
		X"7e", X"7a", X"75", X"71", X"6c", X"6a", X"70", X"7d", X"89", X"8e", X"92", X"8d", X"85", X"83", X"7e", X"7b", 
		X"74", X"71", X"6e", X"70", X"7b", X"84", X"8c", X"91", X"8f", X"89", X"85", X"83", X"81", X"7f", X"7e", X"7b", 
		X"76", X"79", X"83", X"8d", X"95", X"9a", X"95", X"8d", X"88", X"82", X"7e", X"7e", X"7f", X"7d", X"7d", X"7d", 
		X"78", X"72", X"6f", X"6d", X"6c", X"72", X"7f", X"8c", X"90", X"96", X"91", X"88", X"85", X"7f", X"7b", X"74", 
		X"72", X"70", X"70", X"7b", X"84", X"8c", X"91", X"91", X"8b", X"86", X"83", X"80", X"7e", X"7d", X"7a", X"75", 
		X"78", X"81", X"8b", X"95", X"9b", X"97", X"8e", X"88", X"81", X"7d", X"7c", X"7d", X"7b", X"7c", X"7d", X"79", 
		X"74", X"72", X"6f", X"6d", X"72", X"7e", X"8b", X"90", X"95", X"91", X"88", X"84", X"7e", X"7a", X"74", X"72", 
		X"70", X"6f", X"79", X"82", X"8a", X"90", X"90", X"8b", X"85", X"82", X"7e", X"7b", X"7b", X"79", X"75", X"77", 
		X"7e", X"89", X"92", X"99", X"97", X"8f", X"87", X"80", X"7b", X"7a", X"7c", X"7b", X"7c", X"7c", X"79", X"75", 
		X"72", X"71", X"6f", X"71", X"7a", X"87", X"8d", X"93", X"93", X"8b", X"86", X"80", X"7b", X"75", X"72", X"71", 
		X"6f", X"75", X"7e", X"86", X"8d", X"90", X"8e", X"89", X"84", X"7f", X"7b", X"7a", X"79", X"76", X"76", X"7d", 
		X"86", X"8f", X"97", X"98", X"91", X"89", X"81", X"7c", X"7a", X"7d", X"7e", X"7f", X"7f", X"7d", X"78", X"75", 
		X"74", X"71", X"71", X"77", X"83", X"8d", X"93", X"97", X"90", X"89", X"82", X"7c", X"77", X"72", X"72", X"70", 
		X"73", X"7c", X"84", X"8d", X"92", X"93", X"8e", X"87", X"81", X"7b", X"78", X"78", X"76", X"75", X"79", X"82", 
		X"8b", X"94", X"9a", X"97", X"90", X"88", X"80", X"7b", X"7c", X"7d", X"7e", X"7f", X"7f", X"7b", X"77", X"75", 
		X"73", X"72", X"76", X"7f", X"8a", X"90", X"95", X"92", X"8a", X"85", X"7e", X"7a", X"75", X"73", X"72", X"72", 
		X"79", X"81", X"88", X"8e", X"90", X"8d", X"86", X"81", X"7c", X"79", X"78", X"77", X"75", X"77", X"7e", X"87", 
		X"91", X"99", X"99", X"93", X"8a", X"81", X"7b", X"7a", X"7c", X"7e", X"7f", X"7f", X"7e", X"79", X"76", X"75", 
		X"71", X"71", X"76", X"80", X"89", X"8f", X"93", X"8e", X"87", X"81", X"7b", X"77", X"73", X"72", X"71", X"73", 
		X"7a", X"81", X"88", X"8d", X"8e", X"8a", X"84", X"7f", X"7a", X"78", X"78", X"77", X"77", X"7a", X"82", X"8a", 
		X"93", X"99", X"98", X"91", X"88", X"80", X"7a", X"7a", X"7d", X"7f", X"81", X"80", X"7d", X"78", X"75", X"72", 
		X"70", X"72", X"79", X"84", X"8c", X"91", X"93", X"8d", X"88", X"81", X"7b", X"75", X"71", X"70", X"6f", X"74", 
		X"7c", X"83", X"8b", X"8f", X"8f", X"8a", X"85", X"81", X"7c", X"7a", X"79", X"78", X"78", X"7d", X"85", X"8e", 
		X"96", X"9a", X"97", X"8f", X"87", X"7f", X"7b", X"7c", X"7f", X"81", X"82", X"81", X"7c", X"77", X"74", X"71", 
		X"71", X"74", X"7c", X"87", X"8d", X"93", X"93", X"8d", X"87", X"7f", X"7a", X"74", X"71", X"71", X"70", X"76", 
		X"7d", X"86", X"8d", X"90", X"90", X"8a", X"85", X"80", X"7c", X"7a", X"79", X"77", X"78", X"7e", X"86", X"8f", 
		X"97", X"99", X"96", X"8e", X"86", X"7e", X"7a", X"7b", X"7d", X"7f", X"80", X"7f", X"7b", X"77", X"73", X"70", 
		X"70", X"74", X"7d", X"87", X"8d", X"92", X"90", X"8a", X"85", X"7e", X"7a", X"74", X"70", X"6f", X"70", X"76", 
		X"7e", X"87", X"8d", X"90", X"8f", X"8a", X"85", X"80", X"7a", X"78", X"77", X"75", X"77", X"7d", X"85", X"8e", 
		X"95", X"98", X"95", X"8e", X"86", X"7d", X"7a", X"7a", X"7c", X"7e", X"80", X"7f", X"7a", X"75", X"71", X"6d", 
		X"6f", X"73", X"7d", X"88", X"8e", X"92", X"90", X"8b", X"87", X"80", X"7b", X"74", X"70", X"6f", X"6f", X"76", 
		X"7d", X"86", X"8c", X"8f", X"8f", X"8a", X"86", X"81", X"7c", X"7a", X"79", X"77", X"78", X"7d", X"84", X"8c", 
		X"93", X"97", X"95", X"8f", X"88", X"80", X"7c", X"7c", X"7d", X"7f", X"80", X"7e", X"79", X"75", X"72", X"70", 
		X"72", X"77", X"82", X"8c", X"91", X"94", X"91", X"8b", X"85", X"7e", X"79", X"73", X"70", X"6f", X"70", X"77", 
		X"7e", X"87", X"8d", X"90", X"90", X"8b", X"87", X"81", X"7d", X"7b", X"7a", X"78", X"78", X"7c", X"81", X"8a", 
		X"91", X"96", X"95", X"91", X"8a", X"83", X"7f", X"7e", X"7f", X"81", X"81", X"7f", X"7a", X"75", X"71", X"6f", 
		X"71", X"76", X"80", X"8a", X"90", X"93", X"90", X"8a", X"85", X"7e", X"7a", X"74", X"70", X"6f", X"70", X"76", 
		X"7e", X"86", X"8c", X"8f", X"8e", X"8a", X"85", X"80", X"7b", X"79", X"78", X"78", X"78", X"7b", X"80", X"87", 
		X"8f", X"95", X"96", X"93", X"8d", X"85", X"7f", X"7d", X"7d", X"7e", X"7f", X"7d", X"79", X"74", X"70", X"6d", 
		X"6f", X"74", X"7d", X"88", X"8e", X"92", X"91", X"8b", X"85", X"7f", X"7a", X"75", X"71", X"70", X"6e", X"73", 
		X"7b", X"83", X"8a", X"8e", X"8e", X"8a", X"85", X"81", X"7d", X"7c", X"7b", X"7b", X"7a", X"7b", X"7f", X"85", 
		X"8c", X"93", X"96", X"94", X"8e", X"87", X"80", X"7e", X"7d", X"7f", X"80", X"7f", X"7b", X"76", X"71", X"6e", 
		X"6e", X"72", X"7b", X"86", X"8e", X"92", X"92", X"8d", X"88", X"83", X"7e", X"79", X"73", X"70", X"6d", X"70", 
		X"76", X"7f", X"88", X"8e", X"90", X"8e", X"8a", X"86", X"82", X"7f", X"7e", X"7c", X"7a", X"79", X"7b", X"80", 
		X"87", X"90", X"96", X"97", X"93", X"8c", X"85", X"80", X"7e", X"7e", X"7f", X"7f", X"7c", X"77", X"72", X"6e", 
		X"6d", X"71", X"78", X"84", X"8c", X"91", X"93", X"8f", X"8a", X"85", X"80", X"7c", X"75", X"71", X"6e", X"6d", 
		X"73", X"7a", X"84", X"8c", X"90", X"8f", X"8b", X"87", X"83", X"80", X"7e", X"7d", X"7a", X"78", X"79", X"7b", 
		X"82", X"8c", X"93", X"97", X"96", X"90", X"88", X"81", X"7d", X"7c", X"7c", X"7d", X"7c", X"78", X"73", X"6f", 
		X"6c", X"6e", X"74", X"7f", X"89", X"8e", X"91", X"8e", X"8a", X"86", X"82", X"7f", X"79", X"74", X"6f", X"6c", 
		X"6f", X"74", X"7d", X"86", X"8b", X"8d", X"8b", X"88", X"85", X"82", X"81", X"80", X"7e", X"7b", X"79", X"79", 
		X"7d", X"84", X"8d", X"93", X"95", X"92", X"8c", X"85", X"80", X"7d", X"7d", X"7e", X"7d", X"7a", X"75", X"6f", 
		X"6b", X"6b", X"6f", X"79", X"86", X"8d", X"92", X"92", X"8e", X"8a", X"85", X"82", X"7c", X"76", X"71", X"6b", 
		X"6b", X"70", X"78", X"82", X"8a", X"8f", X"8e", X"8c", X"89", X"86", X"85", X"84", X"81", X"7e", X"7a", X"78", 
		X"79", X"7f", X"87", X"8f", X"95", X"95", X"91", X"8a", X"84", X"80", X"7f", X"7f", X"7f", X"7c", X"77", X"71", 
		X"6c", X"69", X"6c", X"75", X"82", X"8d", X"93", X"95", X"90", X"8c", X"87", X"83", X"80", X"7a", X"75", X"6e", 
		X"6b", X"6d", X"72", X"7c", X"85", X"8c", X"8e", X"8d", X"8a", X"87", X"86", X"86", X"85", X"83", X"7f", X"7b", 
		X"78", X"7a", X"81", X"89", X"90", X"93", X"92", X"8c", X"87", X"82", X"7f", X"7f", X"7f", X"7d", X"79", X"72", 
		X"6b", X"67", X"68", X"71", X"7f", X"8a", X"93", X"95", X"90", X"8b", X"86", X"84", X"81", X"7d", X"78", X"70", 
		X"6b", X"69", X"6d", X"76", X"80", X"89", X"8d", X"8d", X"8b", X"87", X"86", X"87", X"87", X"85", X"82", X"7d", 
		X"78", X"78", X"7b", X"82", X"8a", X"90", X"90", X"8d", X"88", X"82", X"7f", X"7e", X"7f", X"7d", X"7a", X"74", 
		X"6b", X"66", X"66", X"6f", X"7c", X"88", X"92", X"94", X"90", X"8c", X"86", X"84", X"82", X"81", X"7c", X"74", 
		X"6e", X"69", X"6b", X"72", X"7b", X"85", X"8b", X"8e", X"8c", X"89", X"88", X"88", X"89", X"8a", X"88", X"82", 
		X"7d", X"79", X"7a", X"7f", X"86", X"8c", X"8f", X"8d", X"89", X"83", X"7f", X"7e", X"7e", X"7e", X"7c", X"76", 
		X"6e", X"68", X"69", X"72", X"7d", X"8a", X"92", X"93", X"90", X"8a", X"85", X"82", X"82", X"82", X"7e", X"79", 
		X"73", X"6d", X"6d", X"71", X"7a", X"82", X"8a", X"8e", X"8c", X"8a", X"88", X"88", X"89", X"8b", X"8a", X"86", 
		X"82", X"7d", X"7c", X"7f", X"84", X"89", X"8c", X"8c", X"88", X"82", X"7f", X"7c", X"7b", X"7b", X"7a", X"75", 
		X"70", X"6e", X"71", X"76", X"81", X"8b", X"8f", X"91", X"8d", X"88", X"83", X"7f", X"80", X"7d", X"7d", X"7a", 
		X"74", X"71", X"6f", X"73", X"78", X"81", X"87", X"8a", X"8b", X"89", X"87", X"86", X"88", X"89", X"88", X"87", 
		X"83", X"80", X"7e", X"7e", X"81", X"84", X"87", X"87", X"85", X"81", X"7d", X"7a", X"78", X"77", X"75", X"72", 
		X"72", X"74", X"77", X"7d", X"85", X"89", X"8c", X"8c", X"89", X"85", X"81", X"7f", X"7c", X"7a", X"7a", X"76", 
		X"75", X"73", X"74", X"77", X"7c", X"82", X"85", X"89", X"8a", X"89", X"88", X"88", X"87", X"86", X"86", X"84", 
		X"82", X"81", X"81", X"81", X"83", X"85", X"85", X"85", X"84", X"80", X"7d", X"7a", X"77", X"75", X"72", X"71", 
		X"74", X"78", X"7e", X"84", X"89", X"8b", X"8c", X"8a", X"87", X"84", X"82", X"80", X"7d", X"7c", X"79", X"77", 
		X"75", X"75", X"77", X"7a", X"7f", X"83", X"86", X"89", X"89", X"89", X"89", X"8a", X"89", X"89", X"88", X"85", 
		X"84", X"82", X"82", X"82", X"84", X"85", X"85", X"84", X"82", X"7f", X"7c", X"79", X"77", X"74", X"73", X"74", 
		X"78", X"7c", X"82", X"88", X"8a", X"8c", X"8a", X"88", X"86", X"83", X"81", X"7e", X"7d", X"7a", X"78", X"77", 
		X"76", X"77", X"78", X"7c", X"80", X"83", X"86", X"88", X"88", X"89", X"89", X"89", X"89", X"88", X"87", X"85", 
		X"84", X"82", X"81", X"81", X"81", X"82", X"82", X"82", X"7f", X"7d", X"7a", X"77", X"74", X"72", X"72", X"76", 
		X"7b", X"80", X"85", X"88", X"89", X"89", X"87", X"85", X"83", X"82", X"7f", X"7d", X"7b", X"79", X"77", X"76", 
		X"76", X"77", X"79", X"7d", X"80", X"83", X"85", X"86", X"87", X"87", X"88", X"88", X"88", X"88", X"86", X"85", 
		X"83", X"81", X"80", X"80", X"81", X"81", X"82", X"80", X"7f", X"7c", X"78", X"75", X"73", X"72", X"74", X"78", 
		X"7d", X"82", X"87", X"88", X"89", X"88", X"86", X"85", X"83", X"82", X"80", X"7f", X"7d", X"7a", X"79", X"77", 
		X"77", X"78", X"7a", X"7d", X"80", X"83", X"85", X"87", X"88", X"88", X"89", X"89", X"89", X"89", X"88", X"87", 
		X"85", X"83", X"82", X"81", X"82", X"82", X"82", X"81", X"80", X"7d", X"79", X"76", X"73", X"73", X"75", X"7a", 
		X"7f", X"85", X"89", X"8a", X"8a", X"88", X"86", X"84", X"83", X"83", X"81", X"80", X"7e", X"7c", X"7a", X"78", 
		X"78", X"78", X"7a", X"7d", X"7f", X"83", X"85", X"86", X"87", X"87", X"88", X"88", X"89", X"89", X"89", X"88", 
		X"86", X"84", X"82", X"81", X"81", X"81", X"82", X"81", X"80", X"7e", X"7a", X"76", X"73", X"72", X"73", X"78", 
		X"7e", X"84", X"88", X"8a", X"89", X"87", X"85", X"83", X"81", X"81", X"81", X"80", X"7f", X"7d", X"7a", X"78", 
		X"76", X"76", X"77", X"7a", X"7c", X"80", X"82", X"84", X"85", X"85", X"86", X"87", X"88", X"89", X"89", X"89", 
		X"87", X"85", X"82", X"80", X"7f", X"7f", X"7f", X"80", X"80", X"7f", X"7c", X"78", X"73", X"71", X"71", X"74", 
		X"7a", X"80", X"86", X"89", X"8a", X"88", X"85", X"83", X"81", X"80", X"80", X"80", X"81", X"7f", X"7e", X"7b", 
		X"78", X"76", X"76", X"77", X"7a", X"7e", X"81", X"84", X"85", X"86", X"86", X"86", X"87", X"88", X"8a", X"8b", 
		X"8a", X"89", X"86", X"83", X"80", X"7f", X"7f", X"7f", X"81", X"81", X"80", X"7d", X"79", X"75", X"72", X"72", 
		X"75", X"7a", X"80", X"86", X"89", X"8a", X"89", X"86", X"83", X"81", X"81", X"81", X"82", X"83", X"82", X"81", 
		X"7e", X"7a", X"77", X"76", X"76", X"79", X"7d", X"81", X"84", X"87", X"88", X"87", X"87", X"87", X"88", X"8a", 
		X"8c", X"8c", X"8c", X"89", X"86", X"82", X"7f", X"7e", X"7e", X"7f", X"81", X"81", X"7f", X"7c", X"78", X"74", 
		X"72", X"73", X"76", X"7c", X"82", X"87", X"89", X"8a", X"88", X"85", X"82", X"80", X"7f", X"7f", X"81", X"82", 
		X"82", X"80", X"7d", X"7a", X"76", X"75", X"75", X"78", X"7c", X"80", X"84", X"87", X"87", X"87", X"87", X"87", 
		X"87", X"89", X"8a", X"8b", X"8a", X"88", X"84", X"81", X"7e", X"7d", X"7d", X"7d", X"7e", X"7e", X"7d", X"7b", 
		X"78", X"75", X"73", X"73", X"76", X"7a", X"7f", X"84", X"87", X"88", X"87", X"85", X"82", X"80", X"7e", X"7e", 
		X"80", X"81", X"81", X"80", X"7e", X"7b", X"78", X"76", X"75", X"77", X"7a", X"7e", X"82", X"85", X"87", X"88", 
		X"88", X"89", X"89", X"89", X"89", X"89", X"88", X"86", X"84", X"82", X"80", X"7f", X"7e", X"7e", X"7e", X"7e", 
		X"7d", X"7c", X"7a", X"79", X"77", X"76", X"77", X"7a", X"7d", X"81", X"84", X"87", X"87", X"86", X"85", X"82", 
		X"81", X"80", X"80", X"81", X"81", X"81", X"80", X"7f", X"7d", X"7b", X"7a", X"7a", X"7b", X"7d", X"80", X"83", 
		X"86", X"89", X"8a", X"8b", X"8b", X"8a", X"89", X"88", X"87", X"86", X"85", X"84", X"83", X"82", X"80", X"7f", 
		X"7e", X"7e", X"7e", X"7d", X"7d", X"7b", X"7a", X"79", X"78", X"79", X"7a", X"7d", X"80", X"83", X"85", X"86", 
		X"86", X"85", X"83", X"82", X"80", X"80", X"80", X"80", X"80", X"80", X"7f", X"7e", X"7d", X"7c", X"7b", X"7b", 
		X"7c", X"7f", X"82", X"86", X"89", X"8a", X"8b", X"8a", X"89", X"87", X"86", X"85", X"84", X"83", X"83", X"82", 
		X"81", X"80", X"7f", X"7e", X"7d", X"7d", X"7c", X"7b", X"7a", X"7a", X"79", X"79", X"79", X"7a", X"7c", X"7e", 
		X"81", X"82", X"84", X"84", X"83", X"83", X"81", X"80", X"7f", X"7f", X"7f", X"7f", X"80", X"7f", X"7f", X"7d", 
		X"7c", X"7c", X"7c", X"7d", X"7f", X"81", X"84", X"86", X"88", X"89", X"89", X"88", X"87", X"85", X"84", X"82", 
		X"81", X"81", X"81", X"82", X"81", X"81", X"80", X"7f", X"7e", X"7d", X"7c", X"7b", X"7a", X"7a", X"7a", X"7b", 
		X"7c", X"7d", X"7e", X"80", X"81", X"82", X"82", X"83", X"83", X"82", X"82", X"82", X"81", X"81", X"81", X"81", 
		X"81", X"80", X"80", X"7f", X"7f", X"7f", X"7f", X"80", X"81", X"83", X"85", X"87", X"88", X"89", X"88", X"87", 
		X"86", X"84", X"83", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"80", X"7f", X"7e", X"7d", X"7d", X"7c", 
		X"7c", X"7c", X"7c", X"7c", X"7c", X"7d", X"7e", X"7f", X"81", X"82", X"83", X"83", X"84", X"83", X"83", X"82", 
		X"82", X"82", X"82", X"82", X"81", X"81", X"80", X"80", X"7f", X"7f", X"80", X"81", X"82", X"84", X"85", X"86", 
		X"87", X"87", X"86", X"85", X"83", X"82", X"82", X"81", X"81", X"82", X"81", X"81", X"80", X"80", X"7f", X"7e", 
		X"7d", X"7d", X"7c", X"7c", X"7b", X"7b", X"7a", X"7a", X"7b", X"7b", X"7d", X"7e", X"7f", X"81", X"82", X"82", 
		X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"7f", X"7f", X"80", X"81", 
		X"82", X"83", X"84", X"85", X"84", X"84", X"83", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"80", X"80", 
		X"80", X"7f", X"7f", X"7e", X"7e", X"7d", X"7d", X"7c", X"7c", X"7b", X"7b", X"7b", X"7b", X"7c", X"7e", X"7f", 
		X"81", X"82", X"83", X"83", X"82", X"82", X"81", X"81", X"81", X"81", X"82", X"83", X"83", X"83", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"82", X"82", X"82", X"81", X"81", 
		X"81", X"81", X"81", X"82", X"81", X"81", X"81", X"80", X"80", X"7f", X"7f", X"7e", X"7d", X"7d", X"7d", X"7d", 
		X"7e", X"7f", X"80", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"83", X"83", X"83", X"83", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"81", X"81", X"80", X"7f", X"7e", 
		X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7f", X"7f", X"80", X"80", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"80", X"80", X"7f", X"7f", 
		X"80", X"80", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"80", X"80", X"7f", X"7f", X"7f", X"7f", X"7f", X"80", X"80", X"80", X"7f", X"7f", X"7f", 
		X"80", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"83", X"83", X"84", X"84", X"84", X"83", X"83", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"83", X"83", X"83", X"83", X"83", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"80", X"80", X"80", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"80", 
		X"80", X"80", X"81", X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"80", 
		X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", 
		X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", 
		X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", 
		X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", 
		X"7d", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", 
		X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7c", X"7c", X"7c", X"7c", 
		X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", 
		X"7c", X"7c", X"7d", X"7d", X"7d", X"7d", X"7e", X"7e", X"7e", X"7e", X"7e", X"7d", X"7d", X"7d", X"7d", X"7d", 
		X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7e", 
		X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", 
		X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"83", X"83", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", 
		X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", 
		X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"82", 
		X"82", X"82", X"83", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", 
		X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"84", X"83", X"83", X"83", 
		X"83", X"83", X"84", X"84", X"84", X"84", X"84", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"82", 
		X"82", X"82", X"82", X"83", X"83", X"83", X"83", X"83", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"7f", X"7f", X"7f", X"7f", X"80", X"80", X"80", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7d", 
		X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7c", X"7c", X"7c", X"7c", X"7c", 
		X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", 
		X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", 
		X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", 
		X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"79", X"79", X"79", X"79", 
		X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", 
		X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"79", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", 
		X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7a", X"7b", X"7b", 
		X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", 
		X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", X"7b", 
		X"7b", X"7b", X"7b", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", 
		X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", 
		X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", 
		X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", X"7c", 
		X"7c", X"7c", X"7c", X"7c", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", 
		X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7d", X"7e", 
		X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"7f", X"7f", X"7f", X"7f", X"7f", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"81", 
		X"80", X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", 
		X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"81", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", 
		X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"83", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"80", X"80", X"80", X"80", 
		X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", 
		X"80", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", X"81", 
		X"81", X"81", X"81", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", 
		X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82", X"82");
	begin
		if rising_edge(clk25) then
			if(sampleCounter >= 3125) then
				if(currentByte > soundLength) then
					currentByte := 0;
				end if;
				soundByte <= Sound(currentByte);
				currentByte := currentByte + 1;
			end if;
		end if;		
	end process;
end Behavioral;

